module FPMUL(opA_i, opB_i, MUL_o);

endmodule
		